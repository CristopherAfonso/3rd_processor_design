module mult_booth()

  registro4 regA();
  registro4 regM();
  registro3 regQ();
  ffdc q1();

  sum_resta4 alu1();
  uc uc0();

endmodule